module P1_img(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b0111100000_0000111111;
		bitarray[1]  = 20'b0111110000_0011111111;
		bitarray[2]  = 20'b0110111000_0111000011;
		bitarray[3]  = 20'b0110011100_1110000011;
		bitarray[4]  = 20'b0110000000_1110000011;
		bitarray[5]  = 20'b0110000000_1110000011;
		bitarray[6]  = 20'b0110000000_1110000011;
		bitarray[7]  = 20'b0110000000_0111000011;
		bitarray[8]  = 20'b0110000000_0001110011;
		bitarray[9]  = 20'b0110000000_0000111111;

		bitarray[10] = 20'b0110000000_0000001111;
		bitarray[11] = 20'b0110000000_0000000111;
		bitarray[12] = 20'b0110000000_0000000011;
		bitarray[13] = 20'b0110000000_0000000011;
		bitarray[14] = 20'b0110000000_0000000011;
		bitarray[15] = 20'b0110000000_0000000011;
		bitarray[16] = 20'b0110000000_0000000011;
		bitarray[17] = 20'b0110000000_0000000011;
		bitarray[18] = 20'b0110000000_0000000011;
		bitarray[19] = 20'b0110000000_0000000011;
	end
endmodule

module P2_img(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b0011111100_0000111111;
		bitarray[1]  = 20'b0111111110_0011111111;
		bitarray[2]  = 20'b1110000111_0111000011;
		bitarray[3]  = 20'b1100000111_1110000011;
		bitarray[4]  = 20'b0110000000_1110000011;
		bitarray[5]  = 20'b0011000000_1110000011;
		bitarray[6]  = 20'b0011000000_1110000011;
		bitarray[7]  = 20'b0001100000_0111000011;
		bitarray[8]  = 20'b0001100000_0001110011;
		bitarray[9]  = 20'b0000110000_0000111111;

		bitarray[10] = 20'b0000110000_0000001111;
		bitarray[11] = 20'b0000011000_0000000111;
		bitarray[12] = 20'b0000011000_0000000011;
		bitarray[13] = 20'b0000001100_0000000011;
		bitarray[14] = 20'b0000001100_0000000011;
		bitarray[15] = 20'b0000000110_0000000011;
		bitarray[16] = 20'b0000000110_0000000011;
		bitarray[17] = 20'b0000000011_0000000011;
		bitarray[18] = 20'b1111111111_0000000011;
		bitarray[19] = 20'b1111111111_0000000011;
	end
endmodule

module target_img(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b00000001111110000000;
		bitarray[1]  = 20'b00000110000001100000;
		bitarray[2]  = 20'b00011000000000011000;
		bitarray[3]  = 20'b00100001111110000100;
		bitarray[4]  = 20'b00100010000001000100;
		bitarray[5]  = 20'b01000100000000100010;
		bitarray[6]  = 20'b01001000111100010010;
		bitarray[7]  = 20'b10010001000010001001;
		bitarray[8]  = 20'b10010010000001001001;
		bitarray[9]  = 20'b10010010011001001001;
		bitarray[10] = 20'b10010010011001001001;
		bitarray[11] = 20'b10010010000001001001;
		bitarray[12] = 20'b10010001000010001001;
		bitarray[13] = 20'b01001000111100010010;
		bitarray[14] = 20'b01000100000000100010;
		bitarray[15] = 20'b00100010000001000100;
		bitarray[16] = 20'b00100001111110000100;
		bitarray[17] = 20'b00011000000000011000;
		bitarray[18] = 20'b00000110000001100000;
		bitarray[19] = 20'b00000001111110000000;
	end
endmodule

module none20(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b00_0000000000000000_00;
		bitarray[1]  = 20'b00_0000000000000000_00;
		bitarray[2]  = 20'b00_0000000000000000_00;
		bitarray[3]  = 20'b00_0000000000000000_00;
		bitarray[4]  = 20'b00_0000000000000000_00;
		bitarray[5]  = 20'b00_0000000000000000_00;
		bitarray[6]  = 20'b00_0000000000000000_00;
		bitarray[7]  = 20'b00_0000000000000000_00;
		bitarray[8]  = 20'b00_0000000000000000_00;
		bitarray[9]  = 20'b00_0000000000000000_00;
		bitarray[10] = 20'b00_0000000000000000_00;
		bitarray[11] = 20'b00_0000000000000000_00;
		bitarray[12] = 20'b00_0000000000000000_00;
		bitarray[13] = 20'b00_0000000000000000_00;
		bitarray[14] = 20'b00_0000000000000000_00;
		bitarray[15] = 20'b00_0000000000000000_00;
		bitarray[16] = 20'b00_0000000000000000_00;
		bitarray[17] = 20'b00_0000000000000000_00;
		bitarray[18] = 20'b00_0000000000000000_00;
		bitarray[19] = 20'b00_0000000000000000_00;
	end
endmodule

module _0(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b00_0000111111110000_00;
		bitarray[1]  = 20'b00_0001111111111000_00;
		bitarray[2]  = 20'b00_0011100000011100_00;
		bitarray[3]  = 20'b00_0111000000001110_00;
		bitarray[4]  = 20'b00_1110000000000111_00;
		bitarray[5]  = 20'b00_1110000000000111_00;
		bitarray[6]  = 20'b00_1110000000000111_00;
		bitarray[7]  = 20'b00_1110000000000111_00;
		bitarray[8]  = 20'b00_1110000000000111_00;
		bitarray[9]  = 20'b00_1110000000000111_00;
		bitarray[10] = 20'b00_1110000000000111_00;
		bitarray[11] = 20'b00_1110000000000111_00;
		bitarray[12] = 20'b00_1110000000000111_00;
		bitarray[13] = 20'b00_1110000000000111_00;
		bitarray[14] = 20'b00_1110000000000111_00;
		bitarray[15] = 20'b00_1110000000000111_00;
		bitarray[16] = 20'b00_0111000000001110_00;
		bitarray[17] = 20'b00_0011100000011100_00;
		bitarray[18] = 20'b00_0001111111111000_00;
		bitarray[19] = 20'b00_0000111111110000_00;
	end
endmodule

module _1(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b00_0000001111110000_00;
		bitarray[1]  = 20'b00_0000001111111000_00;
		bitarray[2]  = 20'b00_0000001111011100_00;
		bitarray[3]  = 20'b00_0000001111001110_00;
		bitarray[4]  = 20'b00_0000001111000111_00;
		bitarray[5]  = 20'b00_0000001111000000_00;
		bitarray[6]  = 20'b00_0000001111000000_00;
		bitarray[7]  = 20'b00_0000001111000000_00;
		bitarray[8]  = 20'b00_0000001111000000_00;
		bitarray[9]  = 20'b00_0000001111000000_00;
		bitarray[10] = 20'b00_0000001111000000_00;
		bitarray[11] = 20'b00_0000001111000000_00;
		bitarray[12] = 20'b00_0000001111000000_00;
		bitarray[13] = 20'b00_0000001111000000_00;
		bitarray[14] = 20'b00_0000001111000000_00;
		bitarray[15] = 20'b00_0000001111000000_00;
		bitarray[16] = 20'b00_0000001111000000_00;
		bitarray[17] = 20'b00_0000001111000000_00;
		bitarray[18] = 20'b00_1111111111111111_00;
		bitarray[19] = 20'b00_1111111111111111_00;
	end
endmodule

module _2(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b00_0000111111110000_00;
		bitarray[1]  = 20'b00_0001111111111000_00;
		bitarray[2]  = 20'b00_0011100000011100_00;
		bitarray[3]  = 20'b00_0111000000001110_00;
		bitarray[4]  = 20'b00_1110000000000111_00;
		bitarray[5]  = 20'b00_1110000000000000_00;
		bitarray[6]  = 20'b00_0111100000000000_00;
		bitarray[7]  = 20'b00_0011110000000000_00;
		bitarray[8]  = 20'b00_0001111000000000_00;
		bitarray[9]  = 20'b00_0000111100000000_00;
		bitarray[10] = 20'b00_0000011110000000_00;
		bitarray[11] = 20'b00_0000001111000000_00;
		bitarray[12] = 20'b00_0000000111100000_00;
		bitarray[13] = 20'b00_0000000011110000_00;
		bitarray[14] = 20'b00_0000000001111000_00;
		bitarray[15] = 20'b00_0000000000111100_00;
		bitarray[16] = 20'b00_0000000000011110_00;
		bitarray[17] = 20'b00_0000000000001111_00;
		bitarray[18] = 20'b00_1111111111111111_00;
		bitarray[19] = 20'b00_1111111111111111_00;
	end
endmodule

module _3(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b00_0000111111110000_00;
		bitarray[1]  = 20'b00_0001111111111000_00;
		bitarray[2]  = 20'b00_0011100000011100_00;
		bitarray[3]  = 20'b00_0111000000001110_00;
		bitarray[4]  = 20'b00_1110000000000111_00;
		bitarray[5]  = 20'b00_1110000000000000_00;
		bitarray[6]  = 20'b00_0111100000000000_00;
		bitarray[7]  = 20'b00_0001111000000000_00;
		bitarray[8]  = 20'b00_0000011110000000_00;
		bitarray[9]  = 20'b00_0000000111100000_00;
		bitarray[10] = 20'b00_0000000111100000_00;
		bitarray[11] = 20'b00_0000011110000000_00;
		bitarray[12] = 20'b00_0001111000000000_00;
		bitarray[13] = 20'b00_0111100000000000_00;
		bitarray[14] = 20'b00_1110000000000000_00;
		bitarray[15] = 20'b00_1110000000000111_00;
		bitarray[16] = 20'b00_0111000000001110_00;
		bitarray[17] = 20'b00_0011100000011100_00;
		bitarray[18] = 20'b00_0001111111111000_00;
		bitarray[19] = 20'b00_0000111111110000_00;
	end
endmodule

module _4(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b00_0001111000000000_00;
		bitarray[1]  = 20'b00_0000111100000000_00;
		bitarray[2]  = 20'b00_0000011110000000_00;
		bitarray[3]  = 20'b00_0000001111000000_00;
		bitarray[4]  = 20'b00_0001111111100000_00;
		bitarray[5]  = 20'b00_0001111011110000_00;
		bitarray[6]  = 20'b00_0001111001111000_00;
		bitarray[7]  = 20'b00_0001111000111100_00;
		bitarray[8]  = 20'b00_0001111000011110_00;
		bitarray[9]  = 20'b00_0001111000001111_00;
		bitarray[10] = 20'b00_1111111111111111_00;
		bitarray[11] = 20'b00_1111111111111111_00;
		bitarray[12] = 20'b00_1111111111111111_00;
		bitarray[13] = 20'b00_0001111000000000_00;
		bitarray[14] = 20'b00_0001111000000000_00;
		bitarray[15] = 20'b00_0001111000000000_00;
		bitarray[16] = 20'b00_0001111000000000_00;
		bitarray[17] = 20'b00_0001111000000000_00;
		bitarray[18] = 20'b00_0001111000000000_00;
		bitarray[19] = 20'b00_0001111000000000_00;
	end
endmodule

module _5(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b00_1111111111111111_00;
		bitarray[1]  = 20'b00_1111111111111111_00;
		bitarray[2]  = 20'b00_1111111111111111_00;
		bitarray[3]  = 20'b00_0000000000001111_00;
		bitarray[4]  = 20'b00_0000000000001111_00;
		bitarray[5]  = 20'b00_0000000000001111_00;
		bitarray[6]  = 20'b00_0000000000001111_00;
		bitarray[7]  = 20'b00_0000000000001111_00;
		bitarray[8]  = 20'b00_0000000000001111_00;
		bitarray[9]  = 20'b00_0000001111111111_00;
		bitarray[10] = 20'b00_0001111111111111_00;
		bitarray[11] = 20'b00_0111111000000111_00;
		bitarray[12] = 20'b00_1111100000000000_00;
		bitarray[13] = 20'b00_1111000000000000_00;
		bitarray[14] = 20'b00_1111000000000000_00;
		bitarray[15] = 20'b00_1111100000000000_00;
		bitarray[16] = 20'b00_0111110000000000_00;
		bitarray[17] = 20'b00_0011110000000000_00;
		bitarray[18] = 20'b00_0000111111110000_00;
		bitarray[19] = 20'b00_0000000111111111_00;
	end
endmodule

module _6(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b00_0001111000000000_00;
		bitarray[1]  = 20'b00_0000111100000000_00;
		bitarray[2]  = 20'b00_0000011110000000_00;
		bitarray[3]  = 20'b00_0000001111000000_00;
		bitarray[4]  = 20'b00_0000000111100000_00;
		bitarray[5]  = 20'b00_0000000011110000_00;
		bitarray[6]  = 20'b00_0000000001111000_00;
		bitarray[7]  = 20'b00_0000000000111100_00;
		bitarray[8]  = 20'b00_0000011111111110_00;
		bitarray[9]  = 20'b00_0001111111111110_00;
		bitarray[10] = 20'b00_0011110000111111_00;
		bitarray[11] = 20'b00_0111100000011111_00;
		bitarray[12] = 20'b00_1111000000001111_00;
		bitarray[13] = 20'b00_1110000000000111_00;
		bitarray[14] = 20'b00_1110000000000111_00;
		bitarray[15] = 20'b00_1111000000001111_00;
		bitarray[16] = 20'b00_0111100000011110_00;
		bitarray[17] = 20'b00_0011110000111100_00;
		bitarray[18] = 20'b00_0001111111111000_00;
		bitarray[19] = 20'b00_0000011111100000_00;
	end
endmodule

module _7(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b00_1111111111111111_00;
		bitarray[1]  = 20'b00_1111111111111111_00;
		bitarray[2]  = 20'b00_1111111111111111_00;
		bitarray[3]  = 20'b00_1111000000000111_00;
		bitarray[4]  = 20'b00_1110000000000011_00;
		bitarray[5]  = 20'b00_1110000000000000_00;
		bitarray[6]  = 20'b00_1111000000000000_00;
		bitarray[7]  = 20'b00_0111100000000000_00;
		bitarray[8]  = 20'b00_0011110000000000_00;
		bitarray[9]  = 20'b00_0001111000000000_00;
		bitarray[10] = 20'b00_0000111100000000_00;
		bitarray[11] = 20'b00_0000011110000000_00;
		bitarray[12] = 20'b00_0000001111000000_00;
		bitarray[13] = 20'b00_0000000111100000_00;
		bitarray[14] = 20'b00_0000000011110000_00;
		bitarray[15] = 20'b00_0000000001111000_00;
		bitarray[16] = 20'b00_0000000000111100_00;
		bitarray[17] = 20'b00_0000000000011110_00;
		bitarray[18] = 20'b00_0000000000001111_00;
		bitarray[19] = 20'b00_0000000000000111_00;
	end
endmodule

module _8(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b00_0000111111110000_00;
		bitarray[1]  = 20'b00_0011111111111100_00;
		bitarray[2]  = 20'b00_0111100000011110_00;
		bitarray[3]  = 20'b00_1111000000001111_00;
		bitarray[4]  = 20'b00_1111000000001111_00;
		bitarray[5]  = 20'b00_0111100000011110_00;
		bitarray[6]  = 20'b00_0011110000111100_00;
		bitarray[7]  = 20'b00_0001111001111000_00;
		bitarray[8]  = 20'b00_0000111111110000_00;
		bitarray[9]  = 20'b00_0000011111100000_00;
		bitarray[10] = 20'b00_0000011111100000_00;
		bitarray[11] = 20'b00_0000111111110000_00;
		bitarray[12] = 20'b00_0001111001111000_00;
		bitarray[13] = 20'b00_0011110000111100_00;
		bitarray[14] = 20'b00_0111100000011110_00;
		bitarray[15] = 20'b00_1111000000001111_00;
		bitarray[16] = 20'b00_1111000000001111_00;
		bitarray[17] = 20'b00_0111100000011110_00;
		bitarray[18] = 20'b00_0011111111111100_00;
		bitarray[19] = 20'b00_0000111111110000_00;
	end
endmodule

module _9(y, xbits);
	input [4:0] y;
	output [19:0] xbits;
	reg [19:0] bitarray[0:19];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 20'b00_0000011111100000_00;
		bitarray[1]  = 20'b00_0001111111111000_00;
		bitarray[2]  = 20'b00_0011110000111100_00;
		bitarray[3]  = 20'b00_0111100000011110_00;
		bitarray[4]  = 20'b00_1111000000001111_00;
		bitarray[5]  = 20'b00_1110000000000111_00;
		bitarray[6]  = 20'b00_1110000000000111_00;
		bitarray[7]  = 20'b00_1111000000001111_00;
		bitarray[8]  = 20'b00_1111100000011110_00;
		bitarray[9]  = 20'b00_1111110000111100_00;
		bitarray[10] = 20'b00_1111111111111000_00;
		bitarray[11] = 20'b00_0111111111100000_00;
		bitarray[12] = 20'b00_0011110000000000_00;
		bitarray[13] = 20'b00_0001111000000000_00;
		bitarray[14] = 20'b00_0000111100000000_00;
		bitarray[15] = 20'b00_0000011110000000_00;
		bitarray[16] = 20'b00_0000001111000000_00;
		bitarray[17] = 20'b00_0000000111100000_00;
		bitarray[18] = 20'b00_0000000011110000_00;
		bitarray[19] = 20'b00_0000000001111000_00;
	end
endmodule

module _(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_000000000000_000000000000_000;
		bitarray[1]  = 30'b000_000000000000_000000000000_000;
		bitarray[2]  = 30'b000_000000000000_000000000000_000;
		bitarray[3]  = 30'b000_000000000000_000000000000_000;
		bitarray[4]  = 30'b000_000000000000_000000000000_000;
		bitarray[5]  = 30'b000_000000000000_000000000000_000;
		bitarray[6]  = 30'b000_000000000000_000000000000_000;
		bitarray[7]  = 30'b000_000000000000_000000000000_000;
		bitarray[8]  = 30'b000_000000000000_000000000000_000;
		bitarray[9]  = 30'b000_000000000000_000000000000_000;
		bitarray[10] = 30'b000_000000000000_000000000000_000;
		bitarray[11] = 30'b000_000000000000_000000000000_000;
		bitarray[12] = 30'b000_000000000000_000000000000_000;
		bitarray[13] = 30'b000_000000000000_000000000000_000;
		bitarray[14] = 30'b000_000000000000_000000000000_000;
		bitarray[15] = 30'b000_000000000000_000000000000_000;
		bitarray[16] = 30'b000_000000000000_000000000000_000;
		bitarray[17] = 30'b000_000000000000_000000000000_000;
		bitarray[18] = 30'b000_000000000000_000000000000_000;
		bitarray[19] = 30'b000_000000000000_000000000000_000;
		bitarray[20] = 30'b000_000000000000_000000000000_000;
		bitarray[21] = 30'b000_000000000000_000000000000_000;
		bitarray[22] = 30'b000_000000000000_000000000000_000;
		bitarray[23] = 30'b000_000000000000_000000000000_000;
		bitarray[24] = 30'b000_000000000000_000000000000_000;
		bitarray[25] = 30'b000_000000000000_000000000000_000;
		bitarray[26] = 30'b000_000000000000_000000000000_000;
		bitarray[27] = 30'b000_000000000000_000000000000_000;
		bitarray[28] = 30'b000_000000000000_000000000000_000;
		bitarray[29] = 30'b000_000000000000_000000000000_000;
	end
endmodule

module W(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_111000000000_000000000111_000;
		bitarray[1]  = 30'b000_111000000000_000000000111_000;
		bitarray[2]  = 30'b000_111000000000_000000000111_000;
		bitarray[3]  = 30'b000_111000000000_000000000111_000;
		bitarray[4]  = 30'b000_111000000000_000000000111_000;
		bitarray[5]  = 30'b000_011100000000_000000001110_000;
		bitarray[6]  = 30'b000_011100000000_000000001110_000;
		bitarray[7]  = 30'b000_011100000000_000000001110_000;
		bitarray[8]  = 30'b000_011100000000_000000001110_000;
		bitarray[9]  = 30'b000_011100000000_000000001110_000;
		bitarray[10] = 30'b000_001110000000_000000011100_000;
		bitarray[11] = 30'b000_001110000000_000000011100_000;
		bitarray[12] = 30'b000_001110000011_110000011100_000;
		bitarray[13] = 30'b000_001110000011_110000011100_000;
		bitarray[14] = 30'b000_001110000011_110000011100_000;
		bitarray[15] = 30'b000_000111000111_111000111000_000;
		bitarray[16] = 30'b000_000111000111_111000111000_000;
		bitarray[17] = 30'b000_000111000111_111000111000_000;
		bitarray[18] = 30'b000_000111000111_111000111000_000;
		bitarray[19] = 30'b000_000111000111_111000111000_000;
		bitarray[20] = 30'b000_000011101110_011101110000_000;
		bitarray[21] = 30'b000_000011101110_011101110000_000;
		bitarray[22] = 30'b000_000011101110_011101110000_000;
		bitarray[23] = 30'b000_000011101110_011101110000_000;
		bitarray[24] = 30'b000_000011101110_011101110000_000;
		bitarray[25] = 30'b000_000001111000_000111100000_000;
		bitarray[26] = 30'b000_000001111000_000111100000_000;
		bitarray[27] = 30'b000_000001111000_000111100000_000;
		bitarray[28] = 30'b000_000001111000_000111100000_000;
		bitarray[29] = 30'b000_000001111000_000111100000_000;
	end
endmodule

module I(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_000011111111_111111110000_000;
		bitarray[1]  = 30'b000_000011111111_111111110000_000;
		bitarray[2]  = 30'b000_000000001111_111100000000_000;
		bitarray[3]  = 30'b000_000000000111_110000000000_000;
		bitarray[4]  = 30'b000_000000000011_110000000000_000;
		bitarray[5]  = 30'b000_000000000011_110000000000_000;
		bitarray[6]  = 30'b000_000000000011_110000000000_000;
		bitarray[7]  = 30'b000_000000000011_110000000000_000;
		bitarray[8]  = 30'b000_000000000011_110000000000_000;
		bitarray[9]  = 30'b000_000000000011_110000000000_000;
		bitarray[10] = 30'b000_000000000011_110000000000_000;
		bitarray[11] = 30'b000_000000000011_110000000000_000;
		bitarray[12] = 30'b000_000000000011_110000000000_000;
		bitarray[13] = 30'b000_000000000011_110000000000_000;
		bitarray[14] = 30'b000_000000000011_110000000000_000;
		bitarray[15] = 30'b000_000000000011_110000000000_000;
		bitarray[16] = 30'b000_000000000011_110000000000_000;
		bitarray[17] = 30'b000_000000000011_110000000000_000;
		bitarray[18] = 30'b000_000000000011_110000000000_000;
		bitarray[19] = 30'b000_000000000011_110000000000_000;
		bitarray[20] = 30'b000_000000000011_110000000000_000;
		bitarray[21] = 30'b000_000000000011_110000000000_000;
		bitarray[22] = 30'b000_000000000011_110000000000_000;
		bitarray[23] = 30'b000_000000000011_110000000000_000;
		bitarray[24] = 30'b000_000000000011_110000000000_000;
		bitarray[25] = 30'b000_000000000011_110000000000_000;
		bitarray[26] = 30'b000_000000000111_111000000000_000;
		bitarray[27] = 30'b000_000000001111_111100000000_000;
		bitarray[28] = 30'b000_000011111111_111111110000_000;
		bitarray[29] = 30'b000_000011111111_111111110000_000;
	end
endmodule

module N(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_111100000000_000000111111_000;
		bitarray[1]  = 30'b000_111100000000_000001111111_000;
		bitarray[2]  = 30'b000_111100000000_000001111111_000;
		bitarray[3]  = 30'b000_111100000000_000011101111_000;
		bitarray[4]  = 30'b000_111100000000_000011101111_000;
		bitarray[5]  = 30'b000_111100000000_000111001111_000;
		bitarray[6]  = 30'b000_111100000000_000111001111_000;
		bitarray[7]  = 30'b000_111100000000_001110001111_000;
		bitarray[8]  = 30'b000_111100000000_001110001111_000;
		bitarray[9]  = 30'b000_111100000000_011100001111_000;
		bitarray[10] = 30'b000_111100000000_011100001111_000;
		bitarray[11] = 30'b000_111100000000_111000001111_000;
		bitarray[12] = 30'b000_111100000000_111000001111_000;
		bitarray[13] = 30'b000_111100000001_110000001111_000;
		bitarray[14] = 30'b000_111100000001_110000001111_000;
		bitarray[15] = 30'b000_111100000011_100000001111_000;
		bitarray[16] = 30'b000_111100000011_100000001111_000;
		bitarray[17] = 30'b000_111100000111_000000001111_000;
		bitarray[18] = 30'b000_111100000111_000000001111_000;
		bitarray[19] = 30'b000_111100001110_000000001111_000;
		bitarray[20] = 30'b000_111100001110_000000001111_000;
		bitarray[21] = 30'b000_111100011100_000000001111_000;
		bitarray[22] = 30'b000_111100011100_000000001111_000;
		bitarray[23] = 30'b000_111100111000_000000001111_000;
		bitarray[24] = 30'b000_111100111000_000000001111_000;
		bitarray[25] = 30'b000_111101110000_000000001111_000;
		bitarray[26] = 30'b000_111101110000_000000001111_000;
		bitarray[27] = 30'b000_111111100000_000000001111_000;
		bitarray[28] = 30'b000_111111100000_000000001111_000;
		bitarray[29] = 30'b000_111111000000_000000001111_000;
	end
endmodule

module L(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_000000000000_000000011111_000;
		bitarray[1]  = 30'b000_000000000000_000000011111_000;
		bitarray[2]  = 30'b000_000000000000_000000011111_000;
		bitarray[3]  = 30'b000_000000000000_000000011111_000;
		bitarray[4]  = 30'b000_000000000000_000000011111_000;
		bitarray[5]  = 30'b000_000000000000_000000011111_000;
		bitarray[6]  = 30'b000_000000000000_000000011111_000;
		bitarray[7]  = 30'b000_000000000000_000000011111_000;
		bitarray[8]  = 30'b000_000000000000_000000011111_000;
		bitarray[9]  = 30'b000_000000000000_000000011111_000;
		bitarray[10] = 30'b000_000000000000_000000011111_000;
		bitarray[11] = 30'b000_000000000000_000000011111_000;
		bitarray[12] = 30'b000_000000000000_000000011111_000;
		bitarray[13] = 30'b000_000000000000_000000011111_000;
		bitarray[14] = 30'b000_000000000000_000000011111_000;
		bitarray[15] = 30'b000_000000000000_000000011111_000;
		bitarray[16] = 30'b000_000000000000_000000011111_000;
		bitarray[17] = 30'b000_000000000000_000000011111_000;
		bitarray[18] = 30'b000_000000000000_000000011111_000;
		bitarray[19] = 30'b000_000000000000_000000011111_000;
		bitarray[20] = 30'b000_000000000000_000000011111_000;
		bitarray[21] = 30'b000_000000000000_000000011111_000;
		bitarray[22] = 30'b000_000000000000_000000011111_000;
		bitarray[23] = 30'b000_000000000000_000000011111_000;
		bitarray[24] = 30'b000_000000000000_000000011111_000;
		bitarray[25] = 30'b000_000000000000_000000011111_000;
		bitarray[26] = 30'b000_111111111111_111111111111_000;
		bitarray[27] = 30'b000_111111111111_111111111111_000;
		bitarray[28] = 30'b000_111111111111_111111111111_000;
		bitarray[29] = 30'b000_111111111111_111111111111_000;
	end
endmodule

module O(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_000000000111_111000000000_000;
		bitarray[1]  = 30'b000_000000011111_111110000000_000;
		bitarray[2]  = 30'b000_000001111111_111111100000_000;
		bitarray[3]  = 30'b000_000011111111_111111110000_000;
		bitarray[4]  = 30'b000_000111111000_000111111000_000;
		bitarray[5]  = 30'b000_000111100000_000001111000_000;
		bitarray[6]  = 30'b000_001111100000_000001111100_000;
		bitarray[7]  = 30'b000_011111000000_000000111110_000;
		bitarray[8]  = 30'b000_011110000000_000000011110_000;
		bitarray[9]  = 30'b000_011110000000_000000011110_000;
		bitarray[10] = 30'b000_111110000000_000000011111_000;
		bitarray[11] = 30'b000_111100000000_000000001111_000;
		bitarray[12] = 30'b000_111100000000_000000001111_000;
		bitarray[13] = 30'b000_111100000000_000000001111_000;
		bitarray[14] = 30'b000_111100000000_000000001111_000;
		bitarray[15] = 30'b000_111100000000_000000001111_000;
		bitarray[16] = 30'b000_111100000000_000000001111_000;
		bitarray[17] = 30'b000_111100000000_000000001111_000;
		bitarray[18] = 30'b000_111100000000_000000001111_000;
		bitarray[19] = 30'b000_111110000000_000000011111_000;
		bitarray[20] = 30'b000_011110000000_000000011110_000;
		bitarray[21] = 30'b000_011110000000_000000011110_000;
		bitarray[22] = 30'b000_011111000000_000000111110_000;
		bitarray[23] = 30'b000_001111100000_000001111100_000;
		bitarray[24] = 30'b000_000111100000_000001111000_000;
		bitarray[25] = 30'b000_000111111000_000111111000_000;
		bitarray[26] = 30'b000_000011111111_111111110000_000;
		bitarray[27] = 30'b000_000001111111_111111100000_000;
		bitarray[28] = 30'b000_000000011111_111110000000_000;
		bitarray[29] = 30'b000_000000000111_111000000000_000;
	end
endmodule

module S(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_000001111111111111100000_000;
		bitarray[1]  = 30'b000_000111111111111111111100_000;
		bitarray[2]  = 30'b000_011111111000000011111110_000;
		bitarray[3]  = 30'b000_111110000000000000011111_000;
		bitarray[4]  = 30'b000_111100000000000000011111_000;
		bitarray[5]  = 30'b000_111000000000000000001110_000;
		bitarray[6]  = 30'b000_000000000000000000011110_000;
		bitarray[7]  = 30'b000_000000000000000000111100_000;
		bitarray[8]  = 30'b000_000000000000000001111000_000;
		bitarray[9]  = 30'b000_000000000000000011110000_000;
		bitarray[10] = 30'b000_000000000000000111100000_000;
		bitarray[11] = 30'b000_000000000000001111000000_000;
		bitarray[12] = 30'b000_000000000000011110000000_000;
		bitarray[13] = 30'b000_000000000000111100000000_000;
		bitarray[14] = 30'b000_000000000001111000000000_000;
		bitarray[15] = 30'b000_000000000011110000000000_000;
		bitarray[16] = 30'b000_000000001111000000000000_000;
		bitarray[17] = 30'b000_000000011110000000000000_000;
		bitarray[18] = 30'b000_000000111100000000000000_000;
		bitarray[19] = 30'b000_000001111000000000000000_000;
		bitarray[20] = 30'b000_000011110000000000000000_000;
		bitarray[21] = 30'b000_000111100000000000000000_000;
		bitarray[22] = 30'b000_001111000000000000000111_000;
		bitarray[23] = 30'b000_111110000000000000001111_000;
		bitarray[24] = 30'b000_111100000000000000001111_000;
		bitarray[25] = 30'b000_111000000000000000001111_000;
		bitarray[26] = 30'b000_111100000000000000111111_000;
		bitarray[27] = 30'b000_011111110000000011111100_000;
		bitarray[28] = 30'b000_000111111111111111111000_000;
		bitarray[29] = 30'b000_000001111111111111110000_000;
	end
endmodule

module E(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_111111111111_111111111111_000;
		bitarray[1]  = 30'b000_111111111111_111111111111_000;
		bitarray[2]  = 30'b000_111111111111_111111111111_000;
		bitarray[3]  = 30'b000_000000000000_000000000111_000;
		bitarray[4]  = 30'b000_000000000000_000000000111_000;
		bitarray[5]  = 30'b000_000000000000_000000000111_000;
		bitarray[6]  = 30'b000_000000000000_000000000111_000;
		bitarray[7]  = 30'b000_000000000000_000000000111_000;
		bitarray[8]  = 30'b000_000000000000_000000000111_000;
		bitarray[9]  = 30'b000_000000000000_000000000111_000;
		bitarray[10] = 30'b000_000000000000_000000000111_000;
		bitarray[11] = 30'b000_000000000000_000000000111_000;
		bitarray[12] = 30'b000_000000000000_000000000111_000;
		bitarray[13] = 30'b000_000000000000_000000000111_000;
		bitarray[14] = 30'b000_000011111111_111111111111_000;
		bitarray[15] = 30'b000_000011111111_111111111111_000;
		bitarray[16] = 30'b000_000011111111_111111111111_000;
		bitarray[17] = 30'b000_000000000000_000000000111_000;
		bitarray[18] = 30'b000_000000000000_000000000111_000;
		bitarray[19] = 30'b000_000000000000_000000000111_000;
		bitarray[20] = 30'b000_000000000000_000000000111_000;
		bitarray[21] = 30'b000_000000000000_000000000111_000;
		bitarray[22] = 30'b000_000000000000_000000000111_000;
		bitarray[23] = 30'b000_000000000000_000000000111_000;
		bitarray[24] = 30'b000_000000000000_000000000111_000;
		bitarray[25] = 30'b000_000000000000_000000000111_000;
		bitarray[26] = 30'b000_000000000000_000000000111_000;
		bitarray[27] = 30'b000_111111111111_111111111111_000;
		bitarray[28] = 30'b000_111111111111_111111111111_000;
		bitarray[29] = 30'b000_111111111111_111111111111_000;
	end
endmodule

module Y(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_111100000000_000000001111_000;
		bitarray[1]  = 30'b000_111100000000_000000001111_000;
		bitarray[2]  = 30'b000_001111000000_000000111100_000;
		bitarray[3]  = 30'b000_001111000000_000000111100_000;
		bitarray[4]  = 30'b000_000011110000_000011110000_000;
		bitarray[5]  = 30'b000_000011110000_000011110000_000;
		bitarray[6]  = 30'b000_000000111100_001111000000_000;
		bitarray[7]  = 30'b000_000000111100_001111000000_000;
		bitarray[8]  = 30'b000_000000001111_111100000000_000;
		bitarray[9]  = 30'b000_000000001111_111100000000_000;
		bitarray[10] = 30'b000_000000000011_110000000000_000;
		bitarray[11] = 30'b000_000000000011_110000000000_000;
		bitarray[12] = 30'b000_000000000011_110000000000_000;
		bitarray[13] = 30'b000_000000000011_110000000000_000;
		bitarray[14] = 30'b000_000000000011_110000000000_000;
		bitarray[15] = 30'b000_000000000011_110000000000_000;
		bitarray[16] = 30'b000_000000000011_110000000000_000;
		bitarray[17] = 30'b000_000000000011_110000000000_000;
		bitarray[18] = 30'b000_000000000011_110000000000_000;
		bitarray[19] = 30'b000_000000000011_110000000000_000;
		bitarray[20] = 30'b000_000000000011_110000000000_000;
		bitarray[21] = 30'b000_000000000011_110000000000_000;
		bitarray[22] = 30'b000_000000000011_110000000000_000;
		bitarray[23] = 30'b000_000000000011_110000000000_000;
		bitarray[24] = 30'b000_000000000011_110000000000_000;
		bitarray[25] = 30'b000_000000000011_110000000000_000;
		bitarray[26] = 30'b000_000000000011_110000000000_000;
		bitarray[27] = 30'b000_000000000011_110000000000_000;
		bitarray[28] = 30'b000_000000000011_110000000000_000;
		bitarray[29] = 30'b000_000000000010_110000000000_000;
	end
endmodule

module U(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_111100000000_000000001111_000;
		bitarray[1]  = 30'b000_111100000000_000000001111_000;
		bitarray[2]  = 30'b000_111100000000_000000001111_000;
		bitarray[3]  = 30'b000_111100000000_000000001111_000;
		bitarray[4]  = 30'b000_111100000000_000000001111_000;
		bitarray[5]  = 30'b000_111100000000_000000001111_000;
		bitarray[6]  = 30'b000_111100000000_000000001111_000;
		bitarray[7]  = 30'b000_111100000000_000000001111_000;
		bitarray[8]  = 30'b000_111100000000_000000001111_000;
		bitarray[9]  = 30'b000_111100000000_000000001111_000;
		bitarray[10] = 30'b000_111100000000_000000001111_000;
		bitarray[11] = 30'b000_111100000000_000000001111_000;
		bitarray[12] = 30'b000_111100000000_000000001111_000;
		bitarray[13] = 30'b000_111100000000_000000001111_000;
		bitarray[14] = 30'b000_111100000000_000000001111_000;
		bitarray[15] = 30'b000_111100000000_000000001111_000;
		bitarray[16] = 30'b000_111100000000_000000001111_000;
		bitarray[17] = 30'b000_111100000000_000000001111_000;
		bitarray[18] = 30'b000_111100000000_000000001111_000;
		bitarray[19] = 30'b000_111100000000_000000001111_000;
		bitarray[20] = 30'b000_111100000000_000000001111_000;
		bitarray[21] = 30'b000_111100000000_000000001111_000;
		bitarray[22] = 30'b000_111100000000_000000001111_000;
		bitarray[23] = 30'b000_111100000000_000000001111_000;
		bitarray[24] = 30'b000_111100000000_000000001111_000;
		bitarray[25] = 30'b000_111110000000_000000011111_000;
		bitarray[26] = 30'b000_011111110000_000011111110_000;
		bitarray[27] = 30'b000_000111111111_111111111000_000;
		bitarray[28] = 30'b000_000001111111_111111100000_000;
		bitarray[29] = 30'b000_000000011111_111110000000_000;
	end
endmodule

module B(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_000000011111_111111111111_000;
		bitarray[1]  = 30'b000_000000111111_111111111111_000;
		bitarray[2]  = 30'b000_000001111111_111111111111_000;
		bitarray[3]  = 30'b000_000111100000_000000001111_000;
		bitarray[4]  = 30'b000_001111000000_000000001111_000;
		bitarray[5]  = 30'b000_011110000000_000000001111_000;
		bitarray[6]  = 30'b000_111100000000_000000001111_000;
		bitarray[7]  = 30'b000_111100000000_000000001111_000;
		bitarray[8]  = 30'b000_111100000000_000000001111_000;
		bitarray[9]  = 30'b000_011110000000_000000001111_000;
		bitarray[10] = 30'b000_001111000000_000000001111_000;
		bitarray[11] = 30'b000_000111100000_000000001111_000;
		bitarray[12] = 30'b000_000011110000_000000001111_000;
		bitarray[13] = 30'b000_000001111100_000000001111_000;
		bitarray[14] = 30'b000_000000011111_111111111111_000;
		bitarray[15] = 30'b000_000000011111_111111111111_000;
		bitarray[16] = 30'b000_000001111100_000000001111_000;
		bitarray[17] = 30'b000_000011110000_000000001111_000;
		bitarray[18] = 30'b000_000111100000_000000001111_000;
		bitarray[19] = 30'b000_001111000000_000000001111_000;
		bitarray[20] = 30'b000_011110000000_000000001111_000;
		bitarray[21] = 30'b000_111100000000_000000001111_000;
		bitarray[22] = 30'b000_111100000000_000000001111_000;
		bitarray[23] = 30'b000_111100000000_000000001111_000;
		bitarray[24] = 30'b000_011110000000_000000001111_000;
		bitarray[25] = 30'b000_001111000000_000000001111_000;
		bitarray[26] = 30'b000_000111100000_000000001111_000;
		bitarray[27] = 30'b000_000011111111_111111111111_000;
		bitarray[28] = 30'b000_000001111111_111111111111_000;
		bitarray[29] = 30'b000_000000111111_111111111111_000;
	end
endmodule

module A(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_000000000111_111000000000_000;
		bitarray[1]  = 30'b000_000000001111_111100000000_000;
		bitarray[2]  = 30'b000_000000001111_111100000000_000;
		bitarray[3]  = 30'b000_000000011110_011110000000_000;
		bitarray[4]  = 30'b000_000000011110_011110000000_000;
		bitarray[5]  = 30'b000_000000111100_001111000000_000;
		bitarray[6]  = 30'b000_000000111100_001111000000_000;
		bitarray[7]  = 30'b000_000001111000_000111100000_000;
		bitarray[8]  = 30'b000_000001111000_000111100000_000;
		bitarray[9]  = 30'b000_000011110000_000011110000_000;
		bitarray[10] = 30'b000_000011110000_000011110000_000;
		bitarray[11] = 30'b000_000111100000_000001111000_000;
		bitarray[12] = 30'b000_000111100000_000001111000_000;
		bitarray[13] = 30'b000_001111000000_000000111100_000;
		bitarray[14] = 30'b000_001111000000_000000111100_000;
		bitarray[15] = 30'b000_111100000000_000000001111_000;
		bitarray[16] = 30'b000_111100000000_000000001111_000;
		bitarray[17] = 30'b000_111100000000_000000001111_000;
		bitarray[18] = 30'b000_111100000000_000000001111_000;
		bitarray[19] = 30'b000_111111111111_111111111111_000;
		bitarray[20] = 30'b000_111111111111_111111111111_000;
		bitarray[21] = 30'b000_111111111111_111111111111_000;
		bitarray[22] = 30'b000_111111111111_111111111111_000;
		bitarray[23] = 30'b000_111100000000_000000001111_000;
		bitarray[24] = 30'b000_111100000000_000000001111_000;
		bitarray[25] = 30'b000_111100000000_000000001111_000;
		bitarray[26] = 30'b000_111100000000_000000001111_000;
		bitarray[27] = 30'b000_111100000000_000000001111_000;
		bitarray[28] = 30'b000_111100000000_000000001111_000;
		bitarray[29] = 30'b000_111100000000_000000001111_000;
	end
endmodule

module P(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_000001111111_111111111111_000;
		bitarray[1]  = 30'b000_000011111111_111111111111_000;
		bitarray[2]  = 30'b000_000111111111_111111111111_000;
		bitarray[3]  = 30'b000_001111000000_000000001111_000;
		bitarray[4]  = 30'b000_011110000000_000000001111_000;
		bitarray[5]  = 30'b000_011110000000_000000001111_000;
		bitarray[6]  = 30'b000_111100000000_000000001111_000;
		bitarray[7]  = 30'b000_111100000000_000000001111_000;
		bitarray[8]  = 30'b000_111100000000_000000001111_000;
		bitarray[9]  = 30'b000_011110000000_000000001111_000;
		bitarray[10] = 30'b000_011110000000_000000001111_000;
		bitarray[11] = 30'b000_001111000000_000000001111_000;
		bitarray[12] = 30'b000_000111111111_111111111111_000;
		bitarray[13] = 30'b000_000011111111_111111111111_000;
		bitarray[14] = 30'b000_000001111111_111111111111_000;
		bitarray[15] = 30'b000_000000000000_000000001111_000;
		bitarray[16] = 30'b000_000000000000_000000001111_000;
		bitarray[17] = 30'b000_000000000000_000000001111_000;
		bitarray[18] = 30'b000_000000000000_000000001111_000;
		bitarray[19] = 30'b000_000000000000_000000001111_000;
		bitarray[20] = 30'b000_000000000000_000000001111_000;
		bitarray[21] = 30'b000_000000000000_000000001111_000;
		bitarray[22] = 30'b000_000000000000_000000001111_000;
		bitarray[23] = 30'b000_000000000000_000000001111_000;
		bitarray[24] = 30'b000_000000000000_000000001111_000;
		bitarray[25] = 30'b000_000000000000_000000001111_000;
		bitarray[26] = 30'b000_000000000000_000000001111_000;
		bitarray[27] = 30'b000_000000000000_000000001111_000;
		bitarray[28] = 30'b000_000000000000_000000001111_000;
		bitarray[29] = 30'b000_000000000000_000000001111_000;
	end
endmodule

module R(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_000001111111_111111111111_000;
		bitarray[1]  = 30'b000_000011111111_111111111111_000;
		bitarray[2]  = 30'b000_000111111111_111111111111_000;
		bitarray[3]  = 30'b000_001111000000_000000001111_000;
		bitarray[4]  = 30'b000_011110000000_000000001111_000;
		bitarray[5]  = 30'b000_011110000000_000000001111_000;
		bitarray[6]  = 30'b000_111100000000_000000001111_000;
		bitarray[7]  = 30'b000_111100000000_000000001111_000;
		bitarray[8]  = 30'b000_111100000000_000000001111_000;
		bitarray[9]  = 30'b000_011110000000_000000001111_000;
		bitarray[10] = 30'b000_011110000000_000000001111_000;
		bitarray[11] = 30'b000_001111000000_000000001111_000;
		bitarray[12] = 30'b000_000111111111_111111111111_000;
		bitarray[13] = 30'b000_000011111111_111111111111_000;
		bitarray[14] = 30'b000_000001111111_111111111111_000;
		bitarray[15] = 30'b000_000000000000_001111001111_000;
		bitarray[16] = 30'b000_000000000000_011110001111_000;
		bitarray[17] = 30'b000_000000000000_111100001111_000;
		bitarray[18] = 30'b000_000000000001_111000001111_000;
		bitarray[19] = 30'b000_000000000011_110000001111_000;
		bitarray[20] = 30'b000_000000000111_100000001111_000;
		bitarray[21] = 30'b000_000000001111_000000001111_000;
		bitarray[22] = 30'b000_000000011110_000000001111_000;
		bitarray[23] = 30'b000_000000111100_000000001111_000;
		bitarray[24] = 30'b000_000001111000_000000001111_000;
		bitarray[25] = 30'b000_000011110000_000000001111_000;
		bitarray[26] = 30'b000_000111100000_000000001111_000;
		bitarray[27] = 30'b000_001111000000_000000001111_000;
		bitarray[28] = 30'b000_011110000000_000000001111_000;
		bitarray[29] = 30'b000_111100000000_000000001111_000;
	end
endmodule

module C(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_000000001111_111100000000_000;
		bitarray[1]  = 30'b000_000000111111_111111000000_000;
		bitarray[2]  = 30'b000_000001111111_111111100000_000;
		bitarray[3]  = 30'b000_000111100000_000001111000_000;
		bitarray[4]  = 30'b000_001111000000_000000111100_000;
		bitarray[5]  = 30'b000_011110000000_000000011110_000;
		bitarray[6]  = 30'b000_111100000000_000000001111_000;
		bitarray[7]  = 30'b000_111100000000_000000001111_000;
		bitarray[8]  = 30'b000_000000000000_000000001111_000;
		bitarray[9]  = 30'b000_000000000000_000000001111_000;
		bitarray[10] = 30'b000_000000000000_000000001111_000;
		bitarray[11] = 30'b000_000000000000_000000001111_000;
		bitarray[12] = 30'b000_000000000000_000000001111_000;
		bitarray[13] = 30'b000_000000000000_000000001111_000;
		bitarray[14] = 30'b000_000000000000_000000001111_000;

		bitarray[15] = 30'b000_000000000000_000000001111_000;
		bitarray[16] = 30'b000_000000000000_000000001111_000;
		bitarray[17] = 30'b000_000000000000_000000001111_000;
		bitarray[18] = 30'b000_000000000000_000000001111_000;
		bitarray[19] = 30'b000_000000000000_000000001111_000;
		bitarray[20] = 30'b000_000000000000_000000001111_000;
		bitarray[21] = 30'b000_000000000000_000000001111_000;
		bitarray[22] = 30'b000_111100000000_000000001111_000;
		bitarray[23] = 30'b000_111100000000_000000001111_000;
		bitarray[24] = 30'b000_011110000000_000000011110_000;
		bitarray[25] = 30'b000_001111000000_000000111100_000;
		bitarray[26] = 30'b000_000111100000_000001111000_000;
		bitarray[27] = 30'b000_000001111111_111111100000_000;
		bitarray[28] = 30'b000_000000111111_111111000000_000;
		bitarray[29] = 30'b000_000000001111_111100000000_000;
	end
endmodule

module G(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_000000001111_111100000000_000;
		bitarray[1]  = 30'b000_000000111111_111111000000_000;
		bitarray[2]  = 30'b000_000001111111_111111100000_000;
		bitarray[3]  = 30'b000_000111100000_000001111000_000;
		bitarray[4]  = 30'b000_001111000000_000000111100_000;
		bitarray[5]  = 30'b000_011110000000_000000011110_000;
		bitarray[6]  = 30'b000_111100000000_000000001111_000;
		bitarray[7]  = 30'b000_111100000000_000000001111_000;
		bitarray[8]  = 30'b000_000000000000_000000001111_000;
		bitarray[9]  = 30'b000_000000000000_000000001111_000;
		bitarray[10] = 30'b000_000000000000_000000001111_000;
		bitarray[11] = 30'b000_000000000000_000000001111_000;
		bitarray[12] = 30'b000_000000000000_000000001111_000;
		bitarray[13] = 30'b000_000000000000_000000001111_000;
		bitarray[14] = 30'b000_000111111111_000000001111_000;
		bitarray[15] = 30'b000_001111111111_000000001111_000;
		bitarray[16] = 30'b000_011111111111_000000001111_000;
		bitarray[17] = 30'b000_111111111111_000000001111_000;
		bitarray[18] = 30'b000_111110000000_000000001111_000;
		bitarray[19] = 30'b000_111100000000_000000001111_000;
		bitarray[20] = 30'b000_111100000000_000000001111_000;
		bitarray[21] = 30'b000_111100000000_000000001111_000;
		bitarray[22] = 30'b000_111100000000_000000001111_000;
		bitarray[23] = 30'b000_111100000000_000000001111_000;
		bitarray[24] = 30'b000_011110000000_000000011110_000;
		bitarray[25] = 30'b000_001111000000_000000111100_000;
		bitarray[26] = 30'b000_000111100000_000001111000_000;
		bitarray[27] = 30'b000_000001111111_111111100000_000;
		bitarray[28] = 30'b000_000000111111_111111000000_000;
		bitarray[29] = 30'b000_000000001111_111100000000_000;
	end
endmodule

module _1_(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_000000000011111100000000_000;
		bitarray[1]  = 30'b000_000000000011111111000000_000;
		bitarray[2]  = 30'b000_000000000011110011110000_000;
		bitarray[3]  = 30'b000_000000000011110001111000_000;
		bitarray[4]  = 30'b000_000000000011110000111100_000;
		bitarray[5]  = 30'b000_000000000011110000011110_000;
		bitarray[6]  = 30'b000_000000000011110000000000_000;
		bitarray[7]  = 30'b000_000000000011110000000000_000;
		bitarray[8]  = 30'b000_000000000011110000000000_000;
		bitarray[9]  = 30'b000_000000000011110000000000_000;
		bitarray[10] = 30'b000_000000000011110000000000_000;
		bitarray[11] = 30'b000_000000000011110000000000_000;
		bitarray[12] = 30'b000_000000000011110000000000_000;
		bitarray[13] = 30'b000_000000000011110000000000_000;
		bitarray[14] = 30'b000_000000000011110000000000_000;
		bitarray[15] = 30'b000_000000000011110000000000_000;
		bitarray[16] = 30'b000_000000000011110000000000_000;
		bitarray[17] = 30'b000_000000000011110000000000_000;
		bitarray[18] = 30'b000_000000000011110000000000_000;
		bitarray[19] = 30'b000_000000000011110000000000_000;
		bitarray[20] = 30'b000_000000000011110000000000_000;
		bitarray[21] = 30'b000_000000000011110000000000_000;
		bitarray[22] = 30'b000_000000000011110000000000_000;
		bitarray[23] = 30'b000_000000000011110000000000_000;
		bitarray[24] = 30'b000_000000000011110000000000_000;
		bitarray[25] = 30'b000_000000000011110000000000_000;
		bitarray[26] = 30'b000_111111111111111111111111_000;
		bitarray[27] = 30'b000_111111111111111111111111_000;
		bitarray[28] = 30'b000_111111111111111111111111_000;
		bitarray[29] = 30'b000_111111111111111111111111_000;
	end
endmodule

module _2_(y, xbits);
	input [4:0] y;
	output [29:0] xbits;
	reg [29:0] bitarray[0:29];
	assign xbits = bitarray[y];
	initial begin // 20*20
		bitarray[0]  = 30'b000_000001111111111111100000_000;
		bitarray[1]  = 30'b000_000111111111111111111100_000;
		bitarray[2]  = 30'b000_011111111111111111111110_000;
		bitarray[3]  = 30'b000_111111000000000000111111_000;
		bitarray[4]  = 30'b000_111110000000000000011111_000;
		bitarray[5]  = 30'b000_111110000000000000000000_000;
		bitarray[6]  = 30'b000_011110000000000000000000_000;
		bitarray[7]  = 30'b000_001111000000000000000000_000;
		bitarray[8]  = 30'b000_000111100000000000000000_000;
		bitarray[9]  = 30'b000_000011110000000000000000_000;
		bitarray[10] = 30'b000_000001111000000000000000_000;
		bitarray[11] = 30'b000_000000111100000000000000_000;
		bitarray[12] = 30'b000_000000001111000000000000_000;
		bitarray[13] = 30'b000_000000000111100000000000_000;
		bitarray[14] = 30'b000_000000000011110000000000_000;
		bitarray[15] = 30'b000_000000000001111000000000_000;
		bitarray[16] = 30'b000_000000000000111100000000_000;
		bitarray[17] = 30'b000_000000000000011110000000_000;
		bitarray[18] = 30'b000_000000000000001111000000_000;
		bitarray[19] = 30'b000_000000000000000111100000_000;
		bitarray[20] = 30'b000_000000000000000011110000_000;
		bitarray[21] = 30'b000_000000000000000001111000_000;
		bitarray[22] = 30'b000_000000000000000000111100_000;
		bitarray[23] = 30'b000_000000000000000000011110_000;
		bitarray[24] = 30'b000_000000000000000000001111_000;
		bitarray[25] = 30'b000_000000000000000000001111_000;
		bitarray[26] = 30'b000_111111111111111111111111_000;
		bitarray[27] = 30'b000_111111111111111111111111_000;
		bitarray[28] = 30'b000_111111111111111111111111_000;
		bitarray[29] = 30'b000_111111111111111111111111_000;
	end
endmodule